/*
 * Write in SV a simple single cycle CPU
 * Behavioral implementation for register file, memories and ALU but focus on FSM and control path
 */

 module single_port_mem(
     input addr;
     output data;
 );
 endmodule

 module dual_port_mem();
 endmodule

 module ALU();
 endmodule

 module regfile();
 endmodule

 module single_cycle_cpu();
 endmodule
